module Pipeline(
  input wire clk,
  input wire reset
)
