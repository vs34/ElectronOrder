module Loader (
  input wire [31:0] imm,
  input wire [31:0] rd
);
  always
